Contract 
  Declarations
      Subject is Loss to Acme by HU
      Inception is 5 Jun 2014
      Expiration is 4 Jun 2015
      PolicyNum is A5059-3
  Covers 
    100% share of 10M 
  Sublimits
    10000 by Wnd
  